module while_loop ;
  int cnt =6;
  
  initial begin 
    while (cnt > 5 )begin 
      cnt++ ;
    $display ("count = %0d , cnt );
              if (cnt == 15) break ;
              end 
              end 
              
              endmodule 
              
    OUTPUT 
# count = 7
# count = 8
# count = 9
# count = 10
# count = 11
# count = 12
# count = 13
# count = 14
# count = 15
    

    
   
