// An event is triggered at the same time as waiting for the event trigger
module event_example();
  event e1;
  
  task process_A();
    $display("@%0t: Before triggering event e1", $time);
    ->e1;
    $display("@%0t: After triggering event e1", $time);
  endtask
  
  task process_B();
    $display("@%0t: waiting for the event e1", $time);
    @e1;
   //wait(e1.triggered);
    $display("@%0t: event e1 is triggered", $time);
  endtask

  initial begin
    fork
      process_A();
      process_B();
   
    join
  end
endmodule

OUTPUT 
# @0: Before triggering event e1
# @0: After triggering event e1
# @0: waiting for the event e1




  =============================================================================================================================================================================================================

  
module event_example();
  event e1;
  
  task process_A();
    $display("@%0t: Before triggering event e1", $time);
    ->e1;
    $display("@%0t: After triggering event e1", $time);
  endtask
  
  task process_B();
    $display("@%0t: waiting for the event e1", $time);
//     @e1;
    wait(e1.triggered );
    $display("@%0t: event e1 is triggered", $time);
  endtask

  initial begin
    fork
      process_A();
      process_B();
   
    join
  end
endmodule

OUTPUT
# @0: Before triggering event e1
# @0: After triggering event e1
# @0: waiting for the event e1
# @0: event e1 is triggered
