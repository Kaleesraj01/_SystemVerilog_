module Three_D_ex;
  int arr[5][6][7];

  
   initial begin 
     int value = 1 ;
     foreach (arr[i,j,k]) begin
       arr [i][j][k] = value++;
     end 
     
     
     foreach (arr[i,j,k]) begin 
       $display ( "arr[%0d][%0d][%0d]= %0d ", i , j ,k, arr[i][j] [k]);
     end end
endmodule 

/* 0utput 
# KERNEL: arr[0][0][0]= 1 
# KERNEL: arr[0][0][1]= 2 
# KERNEL: arr[0][0][2]= 3 
# KERNEL: arr[0][0][3]= 4 
# KERNEL: arr[0][0][4]= 5 
# KERNEL: arr[0][0][5]= 6 
# KERNEL: arr[0][0][6]= 7 
# KERNEL: arr[0][1][0]= 8 
# KERNEL: arr[0][1][1]= 9 
# KERNEL: arr[0][1][2]= 10 
# KERNEL: arr[0][1][3]= 11 
# KERNEL: arr[0][1][4]= 12 
# KERNEL: arr[0][1][5]= 13 
# KERNEL: arr[0][1][6]= 14 
# KERNEL: arr[0][2][0]= 15 
# KERNEL: arr[0][2][1]= 16 
# KERNEL: arr[0][2][2]= 17 
# KERNEL: arr[0][2][3]= 18 
# KERNEL: arr[0][2][4]= 19 
# KERNEL: arr[0][2][5]= 20 
# KERNEL: arr[0][2][6]= 21 
# KERNEL: arr[0][3][0]= 22 
# KERNEL: arr[0][3][1]= 23 
# KERNEL: arr[0][3][2]= 24 
# KERNEL: arr[0][3][3]= 25 
# KERNEL: arr[0][3][4]= 26 
# KERNEL: arr[0][3][5]= 27 
# KERNEL: arr[0][3][6]= 28 
# KERNEL: arr[0][4][0]= 29 
# KERNEL: arr[0][4][1]= 30 
# KERNEL: arr[0][4][2]= 31 
# KERNEL: arr[0][4][3]= 32 
# KERNEL: arr[0][4][4]= 33 
# KERNEL: arr[0][4][5]= 34 
# KERNEL: arr[0][4][6]= 35 
# KERNEL: arr[0][5][0]= 36 
# KERNEL: arr[0][5][1]= 37 
# KERNEL: arr[0][5][2]= 38 
# KERNEL: arr[0][5][3]= 39 
# KERNEL: arr[0][5][4]= 40 
# KERNEL: arr[0][5][5]= 41 
# KERNEL: arr[0][5][6]= 42 
# KERNEL: arr[1][0][0]= 43 
# KERNEL: arr[1][0][1]= 44 
# KERNEL: arr[1][0][2]= 45 
# KERNEL: arr[1][0][3]= 46 
# KERNEL: arr[1][0][4]= 47 
# KERNEL: arr[1][0][5]= 48 
# KERNEL: arr[1][0][6]= 49 
# KERNEL: arr[1][1][0]= 50 
# KERNEL: arr[1][1][1]= 51 
# KERNEL: arr[1][1][2]= 52 
# KERNEL: arr[1][1][3]= 53 
# KERNEL: arr[1][1][4]= 54 
# KERNEL: arr[1][1][5]= 55 
# KERNEL: arr[1][1][6]= 56 
# KERNEL: arr[1][2][0]= 57 
# KERNEL: arr[1][2][1]= 58 
# KERNEL: arr[1][2][2]= 59 
# KERNEL: arr[1][2][3]= 60 
# KERNEL: arr[1][2][4]= 61 
# KERNEL: arr[1][2][5]= 62 
# KERNEL: arr[1][2][6]= 63 
# KERNEL: arr[1][3][0]= 64 
# KERNEL: arr[1][3][1]= 65 
# KERNEL: arr[1][3][2]= 66 
# KERNEL: arr[1][3][3]= 67 
# KERNEL: arr[1][3][4]= 68 
# KERNEL: arr[1][3][5]= 69 
# KERNEL: arr[1][3][6]= 70 
# KERNEL: arr[1][4][0]= 71 
# KERNEL: arr[1][4][1]= 72 
# KERNEL: arr[1][4][2]= 73 
# KERNEL: arr[1][4][3]= 74 
# KERNEL: arr[1][4][4]= 75 
# KERNEL: arr[1][4][5]= 76 
# KERNEL: arr[1][4][6]= 77 
# KERNEL: arr[1][5][0]= 78 
# KERNEL: arr[1][5][1]= 79 
# KERNEL: arr[1][5][2]= 80 
# KERNEL: arr[1][5][3]= 81 
# KERNEL: arr[1][5][4]= 82 
# KERNEL: arr[1][5][5]= 83 
# KERNEL: arr[1][5][6]= 84 
# KERNEL: arr[2][0][0]= 85 
# KERNEL: arr[2][0][1]= 86 
# KERNEL: arr[2][0][2]= 87 
# KERNEL: arr[2][0][3]= 88 
# KERNEL: arr[2][0][4]= 89 
# KERNEL: arr[2][0][5]= 90 
# KERNEL: arr[2][0][6]= 91 
# KERNEL: arr[2][1][0]= 92 
# KERNEL: arr[2][1][1]= 93 
# KERNEL: arr[2][1][2]= 94 
# KERNEL: arr[2][1][3]= 95 
# KERNEL: arr[2][1][4]= 96 
# KERNEL: arr[2][1][5]= 97 
# KERNEL: arr[2][1][6]= 98 
# KERNEL: arr[2][2][0]= 99 
# KERNEL: arr[2][2][1]= 100 
# KERNEL: arr[2][2][2]= 101 
# KERNEL: arr[2][2][3]= 102 
# KERNEL: arr[2][2][4]= 103 
# KERNEL: arr[2][2][5]= 104 
# KERNEL: arr[2][2][6]= 105 
# KERNEL: arr[2][3][0]= 106 
# KERNEL: arr[2][3][1]= 107 
# KERNEL: arr[2][3][2]= 108 
# KERNEL: arr[2][3][3]= 109 
# KERNEL: arr[2][3][4]= 110 
# KERNEL: arr[2][3][5]= 111 
# KERNEL: arr[2][3][6]= 112 
# KERNEL: arr[2][4][0]= 113 
# KERNEL: arr[2][4][1]= 114 
# KERNEL: arr[2][4][2]= 115 
# KERNEL: arr[2][4][3]= 116 
# KERNEL: arr[2][4][4]= 117 
# KERNEL: arr[2][4][5]= 118 
# KERNEL: arr[2][4][6]= 119 
# KERNEL: arr[2][5][0]= 120 
# KERNEL: arr[2][5][1]= 121 
# KERNEL: arr[2][5][2]= 122 
# KERNEL: arr[2][5][3]= 123 
# KERNEL: arr[2][5][4]= 124 
# KERNEL: arr[2][5][5]= 125 
# KERNEL: arr[2][5][6]= 126 
# KERNEL: arr[3][0][0]= 127 
# KERNEL: arr[3][0][1]= 128 
# KERNEL: arr[3][0][2]= 129 
# KERNEL: arr[3][0][3]= 130 
# KERNEL: arr[3][0][4]= 131 
# KERNEL: arr[3][0][5]= 132 
# KERNEL: arr[3][0][6]= 133 
# KERNEL: arr[3][1][0]= 134 
# KERNEL: arr[3][1][1]= 135 
# KERNEL: arr[3][1][2]= 136 
# KERNEL: arr[3][1][3]= 137 
# KERNEL: arr[3][1][4]= 138 
# KERNEL: arr[3][1][5]= 139 
# KERNEL: arr[3][1][6]= 140 
# KERNEL: arr[3][2][0]= 141 
# KERNEL: arr[3][2][1]= 142 
# KERNEL: arr[3][2][2]= 143 
# KERNEL: arr[3][2][3]= 144 
# KERNEL: arr[3][2][4]= 145 
# KERNEL: arr[3][2][5]= 146 
# KERNEL: arr[3][2][6]= 147 
# KERNEL: arr[3][3][0]= 148 
# KERNEL: arr[3][3][1]= 149 
# KERNEL: arr[3][3][2]= 150 
# KERNEL: arr[3][3][3]= 151 
# KERNEL: arr[3][3][4]= 152 
# KERNEL: arr[3][3][5]= 153 
# KERNEL: arr[3][3][6]= 154 
# KERNEL: arr[3][4][0]= 155 
# KERNEL: arr[3][4][1]= 156 
# KERNEL: arr[3][4][2]= 157 
# KERNEL: arr[3][4][3]= 158 
# KERNEL: arr[3][4][4]= 159 
# KERNEL: arr[3][4][5]= 160 
# KERNEL: arr[3][4][6]= 161 
# KERNEL: arr[3][5][0]= 162 
# KERNEL: arr[3][5][1]= 163 
# KERNEL: arr[3][5][2]= 164 
# KERNEL: arr[3][5][3]= 165 
# KERNEL: arr[3][5][4]= 166 
# KERNEL: arr[3][5][5]= 167 
# KERNEL: arr[3][5][6]= 168 
# KERNEL: arr[4][0][0]= 169 
# KERNEL: arr[4][0][1]= 170 
# KERNEL: arr[4][0][2]= 171 
# KERNEL: arr[4][0][3]= 172 
# KERNEL: arr[4][0][4]= 173 
# KERNEL: arr[4][0][5]= 174 
# KERNEL: arr[4][0][6]= 175 
# KERNEL: arr[4][1][0]= 176 
# KERNEL: arr[4][1][1]= 177 
# KERNEL: arr[4][1][2]= 178 
# KERNEL: arr[4][1][3]= 179 
# KERNEL: arr[4][1][4]= 180 
# KERNEL: arr[4][1][5]= 181 
# KERNEL: arr[4][1][6]= 182 
# KERNEL: arr[4][2][0]= 183 
# KERNEL: arr[4][2][1]= 184 
# KERNEL: arr[4][2][2]= 185 
# KERNEL: arr[4][2][3]= 186 
# KERNEL: arr[4][2][4]= 187 
# KERNEL: arr[4][2][5]= 188 
# KERNEL: arr[4][2][6]= 189 
# KERNEL: arr[4][3][0]= 190 
# KERNEL: arr[4][3][1]= 191 
# KERNEL: arr[4][3][2]= 192 
# KERNEL: arr[4][3][3]= 193 
# KERNEL: arr[4][3][4]= 194 
# KERNEL: arr[4][3][5]= 195 
# KERNEL: arr[4][3][6]= 196 
# KERNEL: arr[4][4][0]= 197 
# KERNEL: arr[4][4][1]= 198 
# KERNEL: arr[4][4][2]= 199 
# KERNEL: arr[4][4][3]= 200 
# KERNEL: arr[4][4][4]= 201 
# KERNEL: arr[4][4][5]= 202 
# KERNEL: arr[4][4][6]= 203 
# KERNEL: arr[4][5][0]= 204 
# KERNEL: arr[4][5][1]= 205 
# KERNEL: arr[4][5][2]= 206 
# KERNEL: arr[4][5][3]= 207 
# KERNEL: arr[4][5][4]= 208 
# KERNEL: arr[4][5][5]= 209 
# KERNEL: arr[4][5][6]= 210 
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
Done
